//////////////************RESET TEST************//////////////
class rst_test;
   task reset_test(ref logic rst);
      #75 rst=1'b1;
    endtask
  endclass
